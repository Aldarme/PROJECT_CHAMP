
library ieee;
use ieee.std_logic_1164.all;

entity ASP_HexDisplay is
	port
	(
		hex_4		: out	std_logic_vector(6 downto 0);
		hex_5		: out	std_logic_vector(6 downto 0);
		inNumb	: in	integer;
		reset		: in std_logic
	);
end entity;

architecture hexArch of ASP_HexDisplay is

begin

 ---------------------------------------------------
 --
 --Don't forget that:
 -- high state is '0'
 -- low	 state is '1'
 --
 ---------------------------------------------------
 display : process (inNumb) is

 begin	
	
	case inNumb is
		
		when 0 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '0';
			hex_4(5) <= '0';
			hex_4(6) <= '1';
			
		when 1 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '1';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '1';
			hex_4(4) <= '1';
			hex_4(5) <= '1';
			hex_4(6) <= '1';
			
		when 2 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '1';
			hex_4(3) <= '0';
			hex_4(4) <= '0';
			hex_4(5) <= '1';
			hex_4(6) <= '0';
			
		when 3 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '1';
			hex_4(5) <= '1';
			hex_4(6) <= '0';
			
		when 4 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '1';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '1';
			hex_4(4) <= '1';
			hex_4(5) <= '0';
			hex_4(6) <= '0';
			
		when 5 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '1';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '1';
			hex_4(5) <= '0';
			hex_4(6) <= '0';
			
		when 6 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '1';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '0';
			hex_4(5) <= '0';
			hex_4(6) <= '0';
			
		when 7 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '1';
			hex_4(4) <= '1';
			hex_4(5) <= '1';
			hex_4(6) <= '1';
			
		when 8 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '0';
			hex_4(5) <= '0';
			hex_4(6) <= '0';
			
		when 9 =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '1';
			hex_4(5) <= '0';
			hex_4(6) <= '0';
			
		when 10 =>
			hex_5(0) <= '1';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '1';
			hex_5(4) <= '1';
			hex_5(5) <= '1';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '0';
			hex_4(5) <= '0';
			hex_4(6) <= '1';
			
		when 11 =>
			hex_5(0) <= '1';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '1';
			hex_5(4) <= '1';
			hex_5(5) <= '1';
			hex_5(6) <= '1';
			
			hex_4(0) <= '1';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '1';
			hex_4(4) <= '1';
			hex_4(5) <= '1';
			hex_4(6) <= '1';			
			
		when 12 =>
			hex_5(0) <= '1';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '1';
			hex_5(4) <= '1';
			hex_5(5) <= '1';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '1';
			hex_4(3) <= '0';
			hex_4(4) <= '0';
			hex_4(5) <= '1';
			hex_4(6) <= '0';
			
		when 13 =>
			hex_5(0) <= '1';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '1';
			hex_5(4) <= '1';
			hex_5(5) <= '1';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '1';
			hex_4(5) <= '1';
			hex_4(6) <= '0';
			
		when 14 =>
			hex_5(0) <= '1';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '1';
			hex_5(4) <= '1';
			hex_5(5) <= '1';
			hex_5(6) <= '1';
			
			hex_4(0) <= '1';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '1';
			hex_4(4) <= '1';
			hex_4(5) <= '0';
			hex_4(6) <= '0';
			
		when 15 =>
			hex_5(0) <= '1';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '1';
			hex_5(4) <= '1';
			hex_5(5) <= '1';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '1';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '1';
			hex_4(5) <= '0';
			hex_4(6) <= '0';			
			
		when others =>
			hex_5(0) <= '0';
			hex_5(1) <= '0';
			hex_5(2) <= '0';
			hex_5(3) <= '0';
			hex_5(4) <= '0';
			hex_5(5) <= '0';
			hex_5(6) <= '1';
			
			hex_4(0) <= '0';
			hex_4(1) <= '0';
			hex_4(2) <= '0';
			hex_4(3) <= '0';
			hex_4(4) <= '0';
			hex_4(5) <= '0';
			hex_4(6) <= '1';
			
			
	end case;
 end process display;

end hexarch;